module FMA (
	input logic [31:0] a_fp,
	input logic [31:0] b_fp,
	input logic [31:0] c_fp,
	
	output logic [31:0] out_fp
);

	logic sign_out, largerMag;
	logic [7:0] exp_out, final_exp;
	logic [23:0] mantissa_a, mantissa_b, mantissa_c, mantissa_mul_norm, final_mantissa;
	logic [47:0] mantissa_mul_out;
	logic [24:0] sum_mants;
	
	int i, offset;
	
	always_comb begin
		mantissa_a = {1'b1, a_fp[22:0]};
		mantissa_b = {1'b1, b_fp[22:0]};
		mantissa_c = {1'b1, c_fp[22:0]};
	
		sign_out = a_fp[31] ^ b_fp[31];
		exp_out = a_fp[30:23] + b_fp[30:23] - 8'h7F;
		mantissa_mul_out = mantissa_a * mantissa_b;
		mantissa_mul_norm = mantissa_mul_out[47:24];
		i = 0;
		
		case (mantissa_mul_norm)
			24'b1??????????????????????? : offset = 1;
			24'b01?????????????????????? : offset = 2;
			24'b001????????????????????? : offset = 3;
			24'b0001???????????????????? : offset = 4;
			24'b00001??????????????????? : offset = 5;
			24'b000001?????????????????? : offset = 6;
			24'b0000001????????????????? : offset = 7;
			24'b00000001???????????????? : offset = 8;
			24'b000000001??????????????? : offset = 9;
			24'b0000000001?????????????? : offset = 10;
			24'b00000000001????????????? : offset = 11;
			24'b000000000001???????????? : offset = 12;
			24'b0000000000001??????????? : offset = 13;
			24'b00000000000001?????????? : offset = 14;
			24'b000000000000001????????? : offset = 15;
			24'b0000000000000001???????? : offset = 16;
			24'b00000000000000001??????? : offset = 17;
			24'b000000000000000001?????? : offset = 18;
			24'b0000000000000000001????? : offset = 19;
			24'b00000000000000000001???? : offset = 20;
			24'b000000000000000000001??? : offset = 21;
			24'b0000000000000000000001?? : offset = 22;
			24'b00000000000000000000001? : offset = 23;
			24'b000000000000000000000001 : offset = 24;
			default: offset = 0;
		endcase;
		mantissa_mul_norm = mantissa_mul_norm << offset;
		exp_out = exp_out - (offset-1);
		
		//num1 = mul_out
		//num2 = c_fp
		// largerMag - 1: c > mul_out, 0: mul_out >= c
		
		if(exp_out < c_fp[30:23]) begin
   			final_exp = c_fp[30:23];
  	 		mantissa_mul_norm = mantissa_mul_norm >> (final_exp - exp_out);
  	 		largerMag = 1'b1;
  	 	end else if (c_fp[30:23] < exp_out) begin
   			final_exp = exp_out;
   			mantissa_c = mantissa_c >> (final_exp - c_fp[30:23]);
   			largerMag = 1'b0;
   		end else begin
   			final_exp = exp_out;
   			if (mantissa_c > mantissa_mul_norm) begin
   				largerMag = 1'b1;
   			end else begin
   				largerMag = 1'b0;
   			end
  	 	end
		
		if ((sign_out == 1'b1) && (c_fp[31] == 1'b1)) begin // two positive so add
   			sum_mants = mantissa_c + mantissa_mul_norm;
   			sign_out = 1'b0;
   		
   			final_mantissa = sum_mants[24:1];
   	   		final_exp = final_exp+1;
  	 	end else if ((sign_out == 1'b1) && (c_fp[31] == 1'b0)) begin
  	 		sum_mants = mantissa_mul_norm - mantissa_c;
  	 		sign_out = largerMag ? 1'b1 : 1'b0;
  	 		
  	 		final_mantissa = sum_mants[23:0];
  	 		final_mantissa = sum_mants[24] ? final_mantissa * -1 : final_mantissa;
  	 	end else if ((sign_out == 1'b0) && (c_fp[31] == 1'b1)) begin
  	 		sum_mants = mantissa_c - mantissa_mul_norm;
  	 		sign_out = largerMag ? 1'b0 : 1'b1;
   		
  	 		final_mantissa = sum_mants[23:0];
  	 		final_mantissa = sum_mants[24] ? final_mantissa * -1 : final_mantissa;
  	 	end else begin
  	 		sum_mants = mantissa_c + mantissa_mul_norm;
  	 		sign_out = 1'b1;
  	 		
  	 		final_mantissa = sum_mants[24:1];
  	 		final_exp = final_exp+1;
  	 	end
  	 	
  	 	case (final_mantissa)
			24'b1??????????????????????? : offset = 1;
			24'b01?????????????????????? : offset = 2;
			24'b001????????????????????? : offset = 3;
			24'b0001???????????????????? : offset = 4;
			24'b00001??????????????????? : offset = 5;
			24'b000001?????????????????? : offset = 6;
			24'b0000001????????????????? : offset = 7;
			24'b00000001???????????????? : offset = 8;
			24'b000000001??????????????? : offset = 9;
			24'b0000000001?????????????? : offset = 10;
			24'b00000000001????????????? : offset = 11;
			24'b000000000001???????????? : offset = 12;
			24'b0000000000001??????????? : offset = 13;
			24'b00000000000001?????????? : offset = 14;
			24'b000000000000001????????? : offset = 15;
			24'b0000000000000001???????? : offset = 16;
			24'b00000000000000001??????? : offset = 17;
			24'b000000000000000001?????? : offset = 18;
			24'b0000000000000000001????? : offset = 19;
			24'b00000000000000000001???? : offset = 20;
			24'b000000000000000000001??? : offset = 21;
			24'b0000000000000000000001?? : offset = 22;
			24'b00000000000000000000001? : offset = 23;
			24'b000000000000000000000001 : offset = 24;
			default: offset = 0;
		endcase;
		final_mantissa = final_mantissa << offset;
		final_exp = final_exp - (offset-1);
		
	end
	
	assign out_fp = {~sign_out, final_exp, final_mantissa[23:1]};

endmodule
