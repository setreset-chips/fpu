module fpu_top (
	input logic [31:0] instruction,
	
	output logic [31:0] fpu_out
);

// Misc.

endmodule
