module fln (
            input logic [31:0] num1,
            output logic [31:0] out1
);


   
   
endmodule
   
