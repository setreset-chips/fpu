/*case (mantissa_mul_norm)
			24'b1??????????????????????? : offset = 1;
			24'b01?????????????????????? : offset = 2;
			24'b001????????????????????? : offset = 3;
			24'b0001???????????????????? : offset = 4;
			24'b00001??????????????????? : offset = 5;
			24'b000001?????????????????? : offset = 6;
			24'b0000001????????????????? : offset = 7;
			24'b00000001???????????????? : offset = 8;
			24'b000000001??????????????? : offset = 9;
			24'b0000000001?????????????? : offset = 10;
			24'b00000000001????????????? : offset = 11;
			24'b000000000001???????????? : offset = 12;
			24'b0000000000001??????????? : offset = 13;
			24'b00000000000001?????????? : offset = 14;
			24'b000000000000001????????? : offset = 15;
			24'b0000000000000001???????? : offset = 16;
			24'b00000000000000001??????? : offset = 17;
			24'b000000000000000001?????? : offset = 18;
			24'b0000000000000000001????? : offset = 19;
			24'b00000000000000000001???? : offset = 20;
			24'b000000000000000000001??? : offset = 21;
			24'b0000000000000000000001?? : offset = 22;
			24'b00000000000000000000001? : offset = 23;
			24'b000000000000000000000001 : offset = 24;
			default: offset = 0;
		endcase;
		mantissa_mul_norm = mantissa_mul_norm << offset;
		exp_out = exp_out - (offset-1);*/
		
/*case (final_mantissa)
			24'b1??????????????????????? : offset = 1;
			24'b01?????????????????????? : offset = 2;
			24'b001????????????????????? : offset = 3;
			24'b0001???????????????????? : offset = 4;
			24'b00001??????????????????? : offset = 5;
			24'b000001?????????????????? : offset = 6;
			24'b0000001????????????????? : offset = 7;
			24'b00000001???????????????? : offset = 8;
			24'b000000001??????????????? : offset = 9;
			24'b0000000001?????????????? : offset = 10;
			24'b00000000001????????????? : offset = 11;
			24'b000000000001???????????? : offset = 12;
			24'b0000000000001??????????? : offset = 13;
			24'b00000000000001?????????? : offset = 14;
			24'b000000000000001????????? : offset = 15;
			24'b0000000000000001???????? : offset = 16;
			24'b00000000000000001??????? : offset = 17;
			24'b000000000000000001?????? : offset = 18;
			24'b0000000000000000001????? : offset = 19;
			24'b00000000000000000001???? : offset = 20;
			24'b000000000000000000001??? : offset = 21;
			24'b0000000000000000000001?? : offset = 22;
			24'b00000000000000000000001? : offset = 23;
			24'b000000000000000000000001 : offset = 24;
			default: offset = 0;
		endcase;
		final_mantissa = final_mantissa << offset;
		final_exp = final_exp - (offset-1);*/
