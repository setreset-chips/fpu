module fexp(
	input logic [31:0] base,
	input logic [31:0] exp,
	
	output logic [31:0] out_num
);

	

endmodule
