module fexp(
	
);
